
`define add_op  7'b0000000  // 7'h0
`define sub_op  7'b0000001  // 7'h1
`define and_op  7'b0000110  // 7'h6
`define or_op   7'b0000010  // 7'h2
`define xor_op  7'b0000100  // 7'h4
`define shl_op  7'b0011000  // 7'h18
`define shr_op  7'b0001000  // 7'h8
`define sra_op  7'h10       // 7'h10
`define blt_op  7'b1100000  // 7'h60
`define bltu_op 7'b1110000
`define bge_op  7'b1111000
`define bgeu_op 7'b1111100
`define beq_op  7'b1111110
`define bne_op  7'b1111111
